----------------------------------------------------------------------------------
-- Order Book PCIe Top - Custom RTL Wrapper
-- Integrates pcie_system (XDMA block design) with pcie_bbo_top
--
-- This wrapper:
--   1. Instantiates pcie_system_wrapper (generated from block design)
--   2. Instantiates pcie_bbo_top (BBO to AXI-Stream converter)
--   3. Connects them together
--   4. Includes test BBO generator for MVP validation
--
-- Target: AX7203 (XC7A200T-2FBG484I)
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity order_book_pcie_top is
    Port (
        -- PCIe interface (directly from FPGA pins)
        pcie_mgt_rxn      : in  STD_LOGIC_VECTOR(3 downto 0);
        pcie_mgt_rxp      : in  STD_LOGIC_VECTOR(3 downto 0);
        pcie_mgt_txn      : out STD_LOGIC_VECTOR(3 downto 0);
        pcie_mgt_txp      : out STD_LOGIC_VECTOR(3 downto 0);

        -- PCIe reference clock (100 MHz differential)
        pcie_refclk_clk_n : in  STD_LOGIC_VECTOR(0 downto 0);
        pcie_refclk_clk_p : in  STD_LOGIC_VECTOR(0 downto 0);

        -- PCIe reset (active low)
        reset_rtl_0       : in  STD_LOGIC;

        -- Status LED
        user_lnk_up       : out STD_LOGIC
    );
end order_book_pcie_top;

architecture Behavioral of order_book_pcie_top is

    -- TEST MODE options (integer to avoid Xilinx boolean synthesis issues):
    -- 0 = Normal BBO mode (pcie_bbo_top with CDC FIFO)
    -- 1 = Simple counter test (continuous incrementing data)
    -- 2 = Direct BBO test (bypass pcie_bbo_top, format BBO packets directly)
    constant TEST_MODE : integer := 2;

    -- Block design wrapper component (generated by Vivado)
    component pcie_system_wrapper is
        Port (
            -- PCIe MGT
            pcie_mgt_rxn      : in  STD_LOGIC_VECTOR(3 downto 0);
            pcie_mgt_rxp      : in  STD_LOGIC_VECTOR(3 downto 0);
            pcie_mgt_txn      : out STD_LOGIC_VECTOR(3 downto 0);
            pcie_mgt_txp      : out STD_LOGIC_VECTOR(3 downto 0);
            -- PCIe clock and reset
            pcie_refclk_clk_n : in  STD_LOGIC_VECTOR(0 downto 0);
            pcie_refclk_clk_p : in  STD_LOGIC_VECTOR(0 downto 0);
            reset_rtl_0       : in  STD_LOGIC;
            -- AXI clock and reset (output from XDMA)
            axi_aclk          : out STD_LOGIC;
            axi_aresetn       : out STD_LOGIC;
            -- S_AXIS_C2H (input from custom logic)
            s_axis_c2h_tdata  : in  STD_LOGIC_VECTOR(63 downto 0);
            s_axis_c2h_tkeep  : in  STD_LOGIC_VECTOR(7 downto 0);
            s_axis_c2h_tlast  : in  STD_LOGIC;
            s_axis_c2h_tready : out STD_LOGIC;
            s_axis_c2h_tvalid : in  STD_LOGIC;
            -- Status
            user_lnk_up       : out STD_LOGIC
        );
    end component;

    -- pcie_bbo_top component (BBO to AXI-Stream converter)
    component pcie_bbo_top is
        Generic (
            C_AXI_DATA_WIDTH      : integer := 64;
            C_AXI_LITE_DATA_WIDTH : integer := 32;
            C_AXI_LITE_ADDR_WIDTH : integer := 6
        );
        Port (
            -- Trading clock domain
            clk_trading    : in  STD_LOGIC;
            rst_trading    : in  STD_LOGIC;
            -- BBO input
            bbo_update     : in  STD_LOGIC;
            bbo_symbol     : in  STD_LOGIC_VECTOR(63 downto 0);
            bbo_bid_price  : in  STD_LOGIC_VECTOR(31 downto 0);
            bbo_bid_size   : in  STD_LOGIC_VECTOR(31 downto 0);
            bbo_ask_price  : in  STD_LOGIC_VECTOR(31 downto 0);
            bbo_ask_size   : in  STD_LOGIC_VECTOR(31 downto 0);
            bbo_spread     : in  STD_LOGIC_VECTOR(31 downto 0);
            -- Timestamps
            ts_t1          : in  STD_LOGIC_VECTOR(31 downto 0);
            ts_t2          : in  STD_LOGIC_VECTOR(31 downto 0);
            ts_t3          : in  STD_LOGIC_VECTOR(31 downto 0);
            ts_t4          : in  STD_LOGIC_VECTOR(31 downto 0);
            -- XDMA clock domain
            axi_aclk       : in  STD_LOGIC;
            axi_aresetn    : in  STD_LOGIC;
            -- AXI-Stream Master (to XDMA C2H)
            m_axis_tdata   : out STD_LOGIC_VECTOR(63 downto 0);
            m_axis_tkeep   : out STD_LOGIC_VECTOR(7 downto 0);
            m_axis_tvalid  : out STD_LOGIC;
            m_axis_tready  : in  STD_LOGIC;
            m_axis_tlast   : out STD_LOGIC;
            -- AXI-Lite Slave (control registers)
            S_AXI_AWADDR   : in  STD_LOGIC_VECTOR(5 downto 0);
            S_AXI_AWVALID  : in  STD_LOGIC;
            S_AXI_AWREADY  : out STD_LOGIC;
            S_AXI_WDATA    : in  STD_LOGIC_VECTOR(31 downto 0);
            S_AXI_WSTRB    : in  STD_LOGIC_VECTOR(3 downto 0);
            S_AXI_WVALID   : in  STD_LOGIC;
            S_AXI_WREADY   : out STD_LOGIC;
            S_AXI_BRESP    : out STD_LOGIC_VECTOR(1 downto 0);
            S_AXI_BVALID   : out STD_LOGIC;
            S_AXI_BREADY   : in  STD_LOGIC;
            S_AXI_ARADDR   : in  STD_LOGIC_VECTOR(5 downto 0);
            S_AXI_ARVALID  : in  STD_LOGIC;
            S_AXI_ARREADY  : out STD_LOGIC;
            S_AXI_RDATA    : out STD_LOGIC_VECTOR(31 downto 0);
            S_AXI_RRESP    : out STD_LOGIC_VECTOR(1 downto 0);
            S_AXI_RVALID   : out STD_LOGIC;
            S_AXI_RREADY   : in  STD_LOGIC;
            -- Status LEDs
            led_link_up    : out STD_LOGIC;
            led_streaming  : out STD_LOGIC;
            led_overflow   : out STD_LOGIC
        );
    end component;

    -- Internal signals
    signal axi_aclk_int       : STD_LOGIC;
    signal axi_aresetn_int    : STD_LOGIC;
    signal rst_trading_int    : STD_LOGIC;

    -- AXI-Stream signals (pcie_bbo_top -> XDMA)
    signal c2h_tdata          : STD_LOGIC_VECTOR(63 downto 0);
    signal c2h_tkeep          : STD_LOGIC_VECTOR(7 downto 0);
    signal c2h_tvalid         : STD_LOGIC;
    signal c2h_tready         : STD_LOGIC;
    signal c2h_tlast          : STD_LOGIC;

    -- Test BBO generator signals
    signal bbo_update_int     : STD_LOGIC;
    signal bbo_timer          : unsigned(23 downto 0) := (others => '0');
    signal bbo_timer_prev     : STD_LOGIC := '0';
    signal bbo_counter        : unsigned(15 downto 0) := (others => '0');

    -- Test BBO data
    constant TEST_SYMBOL      : STD_LOGIC_VECTOR(63 downto 0) := x"544553544141504C"; -- "TESTAAPL"
    signal test_bid_price     : STD_LOGIC_VECTOR(31 downto 0);
    signal test_ask_price     : STD_LOGIC_VECTOR(31 downto 0);
    signal test_timestamp     : STD_LOGIC_VECTOR(31 downto 0);

    -- Simple test pattern signals (for debugging XDMA)
    signal test_counter       : unsigned(63 downto 0) := (others => '0');
    signal test_tdata         : STD_LOGIC_VECTOR(63 downto 0);
    signal test_tvalid        : STD_LOGIC := '0';
    signal test_tlast         : STD_LOGIC := '0';
    signal test_beat_count    : unsigned(2 downto 0) := (others => '0');

    -- Direct BBO test signals (mode 2)
    -- States: 0=IDLE, 1-6=BEAT1-6 (outputs are combinatorial from state)
    signal direct_bbo_state   : integer range 0 to 6 := 0;
    signal direct_bbo_tdata   : STD_LOGIC_VECTOR(63 downto 0) := (others => '0');
    signal direct_bbo_tvalid  : STD_LOGIC := '0';
    signal direct_bbo_tlast   : STD_LOGIC := '0';
    signal direct_bbo_pkt_cnt : unsigned(31 downto 0) := (others => '0');
    signal direct_bbo_timer   : unsigned(19 downto 0) := (others => '0');  -- ~4ms at 250MHz

begin

    -- Trading reset (active high) from axi_aresetn (active low)
    rst_trading_int <= not axi_aresetn_int;

    ---------------------------------------------------------------------------
    -- Block Design Instance (XDMA + clock infrastructure)
    ---------------------------------------------------------------------------
    pcie_system_inst : pcie_system_wrapper
        port map (
            -- PCIe MGT
            pcie_mgt_rxn      => pcie_mgt_rxn,
            pcie_mgt_rxp      => pcie_mgt_rxp,
            pcie_mgt_txn      => pcie_mgt_txn,
            pcie_mgt_txp      => pcie_mgt_txp,
            -- PCIe clock and reset
            pcie_refclk_clk_n => pcie_refclk_clk_n,
            pcie_refclk_clk_p => pcie_refclk_clk_p,
            reset_rtl_0       => reset_rtl_0,
            -- AXI clock and reset
            axi_aclk          => axi_aclk_int,
            axi_aresetn       => axi_aresetn_int,
            -- S_AXIS_C2H (from pcie_bbo_top)
            s_axis_c2h_tdata  => c2h_tdata,
            s_axis_c2h_tkeep  => c2h_tkeep,
            s_axis_c2h_tlast  => c2h_tlast,
            s_axis_c2h_tready => c2h_tready,
            s_axis_c2h_tvalid => c2h_tvalid,
            -- Status
            user_lnk_up       => user_lnk_up
        );

    ---------------------------------------------------------------------------
    -- Test BBO Generator
    -- Generates periodic BBO updates (~250/sec at 250MHz clock)
    ---------------------------------------------------------------------------
    process(axi_aclk_int)
    begin
        if rising_edge(axi_aclk_int) then
            if axi_aresetn_int = '0' then
                bbo_timer <= (others => '0');
                bbo_timer_prev <= '0';
                bbo_counter <= (others => '0');
                bbo_update_int <= '0';
            else
                -- Free-running timer
                bbo_timer <= bbo_timer + 1;
                bbo_timer_prev <= bbo_timer(23);

                -- Generate pulse on MSB edge (~250 updates/sec at 250MHz)
                if bbo_timer(23) = '1' and bbo_timer_prev = '0' then
                    bbo_update_int <= '1';
                    bbo_counter <= bbo_counter + 1;
                else
                    bbo_update_int <= '0';
                end if;
            end if;
        end if;
    end process;

    -- Test prices: Bid = 100.XX, Ask = 101.XX (XX = counter)
    test_bid_price <= x"0064" & std_logic_vector(bbo_counter);
    test_ask_price <= x"0065" & std_logic_vector(bbo_counter);
    test_timestamp <= x"00" & std_logic_vector(bbo_timer);

    ---------------------------------------------------------------------------
    -- pcie_bbo_top Instance (BBO to AXI-Stream converter)
    -- Only instantiated in normal mode (TEST_MODE = 0)
    ---------------------------------------------------------------------------
    gen_bbo_path: if TEST_MODE = 0 generate
        pcie_bbo_inst : pcie_bbo_top
            generic map (
                C_AXI_DATA_WIDTH      => 64,
                C_AXI_LITE_DATA_WIDTH => 32,
                C_AXI_LITE_ADDR_WIDTH => 6
            )
            port map (
                -- Trading clock (use XDMA clock for MVP - no CDC needed)
                clk_trading    => axi_aclk_int,
                rst_trading    => rst_trading_int,
                -- Test BBO data
                bbo_update     => bbo_update_int,
                bbo_symbol     => TEST_SYMBOL,
                bbo_bid_price  => test_bid_price,
                bbo_bid_size   => x"00000064",    -- 100 shares
                bbo_ask_price  => test_ask_price,
                bbo_ask_size   => x"000000C8",    -- 200 shares
                bbo_spread     => x"00010000",    -- 1.0 spread
                -- Timestamps
                ts_t1          => test_timestamp,
                ts_t2          => test_timestamp,
                ts_t3          => test_timestamp,
                ts_t4          => test_timestamp,
                -- XDMA clock domain
                axi_aclk       => axi_aclk_int,
                axi_aresetn    => axi_aresetn_int,
                -- AXI-Stream to XDMA
                m_axis_tdata   => c2h_tdata,
                m_axis_tkeep   => c2h_tkeep,
                m_axis_tvalid  => c2h_tvalid,
                m_axis_tready  => c2h_tready,
                m_axis_tlast   => c2h_tlast,
                -- AXI-Lite (tied off for MVP)
                S_AXI_AWADDR   => (others => '0'),
                S_AXI_AWVALID  => '0',
                S_AXI_AWREADY  => open,
                S_AXI_WDATA    => (others => '0'),
                S_AXI_WSTRB    => (others => '0'),
                S_AXI_WVALID   => '0',
                S_AXI_WREADY   => open,
                S_AXI_BRESP    => open,
                S_AXI_BVALID   => open,
                S_AXI_BREADY   => '0',
                S_AXI_ARADDR   => (others => '0'),
                S_AXI_ARVALID  => '0',
                S_AXI_ARREADY  => open,
                S_AXI_RDATA    => open,
                S_AXI_RRESP    => open,
                S_AXI_RVALID   => open,
                S_AXI_RREADY   => '0',
                -- LEDs (directly from block design for now)
                led_link_up    => open,
                led_streaming  => open,
                led_overflow   => open
            );
    end generate;

    ---------------------------------------------------------------------------
    -- Simple Test Pattern Generator (TEST_MODE = 1)
    -- Generates continuous 64-bit incrementing data with TLAST every 6 beats
    ---------------------------------------------------------------------------
    gen_simple_test: if TEST_MODE = 1 generate
        process(axi_aclk_int)
        begin
            if rising_edge(axi_aclk_int) then
                if axi_aresetn_int = '0' then
                    test_counter <= (others => '0');
                    test_tvalid <= '0';
                    test_tlast <= '0';
                    test_beat_count <= (others => '0');
                else
                    -- Always valid after reset
                    test_tvalid <= '1';

                    -- Increment counter when ready
                    if c2h_tready = '1' then
                        test_counter <= test_counter + 1;
                        test_beat_count <= test_beat_count + 1;

                        -- Assert TLAST every 6 beats (48 bytes = one "packet")
                        if test_beat_count = 5 then
                            test_tlast <= '1';
                            test_beat_count <= (others => '0');
                        else
                            test_tlast <= '0';
                        end if;
                    end if;
                end if;
            end if;
        end process;

        test_tdata <= std_logic_vector(test_counter);

        -- Route test pattern to C2H (override pcie_bbo_top output)
        c2h_tdata  <= test_tdata;
        c2h_tkeep  <= (others => '1');
        c2h_tvalid <= test_tvalid;
        c2h_tlast  <= test_tlast;
    end generate;

    ---------------------------------------------------------------------------
    -- Direct BBO Test Generator (TEST_MODE = 2)
    -- Formats BBO packets directly, bypassing pcie_bbo_top
    -- Sends one 48-byte BBO packet every ~8ms at 125MHz (125 packets/sec)
    --
    -- BYTE ORDER: For AXI-Stream 64-bit to little-endian x86 host:
    --   tdata[7:0]   -> memory byte 0 (first byte in packet)
    --   tdata[63:56] -> memory byte 7
    -- For two 32-bit fields in one 64-bit beat:
    --   First field (lower address) goes in tdata[31:0]
    --   Second field (higher address) goes in tdata[63:32]
    ---------------------------------------------------------------------------
    gen_direct_bbo: if TEST_MODE = 2 generate
        -- Clocked process: only handles state transitions, timer, and packet counter
        -- All AXI-Stream outputs (tdata, tvalid, tlast) are combinatorial from state
        process(axi_aclk_int)
        begin
            if rising_edge(axi_aclk_int) then
                if axi_aresetn_int = '0' then
                    direct_bbo_state <= 0;
                    direct_bbo_pkt_cnt <= (others => '0');
                    direct_bbo_timer <= (others => '0');
                else
                    -- Timer to trigger new packets (~4ms at 250MHz)
                    direct_bbo_timer <= direct_bbo_timer + 1;

                    -- State machine: state transitions only
                    case direct_bbo_state is
                        when 0 =>  -- IDLE - wait for timer
                            if direct_bbo_timer = 0 then
                                direct_bbo_state <= 1;
                            end if;

                        when 1 =>  -- BEAT1: Symbol
                            if c2h_tready = '1' then
                                direct_bbo_state <= 2;
                            end if;

                        when 2 =>  -- BEAT2: BidPrice + BidSize
                            if c2h_tready = '1' then
                                direct_bbo_state <= 3;
                            end if;

                        when 3 =>  -- BEAT3: AskPrice + AskSize
                            if c2h_tready = '1' then
                                direct_bbo_state <= 4;
                            end if;

                        when 4 =>  -- BEAT4: Spread + T1
                            if c2h_tready = '1' then
                                direct_bbo_state <= 5;
                            end if;

                        when 5 =>  -- BEAT5: T2 + T3
                            if c2h_tready = '1' then
                                direct_bbo_state <= 6;
                            end if;

                        when 6 =>  -- BEAT6: T4 + Padding with TLAST
                            if c2h_tready = '1' then
                                direct_bbo_pkt_cnt <= direct_bbo_pkt_cnt + 1;
                                direct_bbo_state <= 0;
                            end if;

                        when others =>
                            direct_bbo_state <= 0;
                    end case;
                end if;
            end if;
        end process;

        -- Combinatorial outputs based on state
        -- All signals change together when state changes, ensuring alignment

        -- tvalid: high for states 1-6 (all beat states)
        direct_bbo_tvalid <= '1' when (direct_bbo_state >= 1 and direct_bbo_state <= 6) else '0';

        -- tlast: high only for state 6 (last beat)
        direct_bbo_tlast <= '1' when direct_bbo_state = 6 else '0';

        -- tdata: select based on state
        with direct_bbo_state select direct_bbo_tdata <=
            -- BEAT1: Symbol "TESTAAPL" (ASCII: 54 45 53 54 41 41 50 4C)
            x"4C50414154534554"                                              when 1,
            -- BEAT2: BidPrice (15000 = $1.50) | BidSize (100)
            x"00000064" & x"00003A98"                                        when 2,
            -- BEAT3: AskPrice (15100 = $1.51) | AskSize (200)
            x"000000C8" & x"00003AFC"                                        when 3,
            -- BEAT4: T1 (pkt_cnt) | Spread (100 = $0.01)
            std_logic_vector(direct_bbo_pkt_cnt) & x"00000064"               when 4,
            -- BEAT5: T3 (pkt_cnt) | T2 (pkt_cnt)
            std_logic_vector(direct_bbo_pkt_cnt) & std_logic_vector(direct_bbo_pkt_cnt) when 5,
            -- BEAT6: Padding (0xDEADBEEF) | T4 (pkt_cnt)
            x"DEADBEEF" & std_logic_vector(direct_bbo_pkt_cnt)               when 6,
            -- Default (IDLE and others)
            x"0000000000000000"                                              when others;

        -- Route direct BBO pattern to C2H
        c2h_tdata  <= direct_bbo_tdata;
        c2h_tkeep  <= (others => '1');
        c2h_tvalid <= direct_bbo_tvalid;
        c2h_tlast  <= direct_bbo_tlast;
    end generate;

end Behavioral;
